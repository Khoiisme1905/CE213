library verilog;
use verilog.vl_types.all;
entity lab_3_mealy_vlg_vec_tst is
end lab_3_mealy_vlg_vec_tst;
