module Instruction_Memory (
    input rst,          // Tin hieu reset
    input [31:0] A,     // Dia chi lenh
    output wire [31:0] RD // Ma lenh doc ra
);
    reg [31:0] mem[0:1023]; // Mang 1024 tu, moi tu 32 bit

    // Khởi tạo bộ nhớ lệnh trực tiếp
    integer i;
    initial begin
        // Khởi tạo tất cả bộ nhớ với giá trị 0
        for (i = 0; i < 1024; i = i + 1) begin
            mem[i] = 32'h00000000;
        end
        
        // Nạp lệnh cho chương trình
        mem[0] = 32'b00000010101000000000001100010011;
        mem[1] = 32'b00000110010000000000001110010011;
        mem[2] = 32'b00000000011001010010000000100011;
        mem[3] = 32'b00000000011101010010001000100011;
        mem[4] = 32'b00000000000001010010111000000011;
        mem[5] = 32'b00000000010001010010111010000011;
        mem[6] = 32'b00000011011100000000111100010011;
        mem[7] = 32'b00000001111001010010010000100011;
        mem[8] = 32'b00000000000001010010111110000011;
        mem[9] = 32'b00000000010001010010001010000011;
        mem[10] = 32'b00000000010111111000111110110011;
        mem[11] = 32'b00000000100001010010001010000011;
        mem[12] = 32'b00000000010111111000111110110011;
        mem[13] = 32'b00000001111101010010011000100011;
    end

    assign RD = (rst == 1'b0) ? {32{1'b0}} : mem[A[31:2]]; // Doc lenh tu dia chi (bo 2 bit thap)
endmodule