library verilog;
use verilog.vl_types.all;
entity lab_3_mealy_vlg_check_tst is
    port(
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_3_mealy_vlg_check_tst;
